module const4 (Y);
	parameter CONST = 0;
	
	output [3:0] Y;
	
	assign Y = CONST; 
	
endmodule