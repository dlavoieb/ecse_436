for j in 0 to NUMBER_OF_SAMPLES-1 loop
    data(j) <= temp(SAMPLES_DATA_LENGTH -5 downto 0) & "0000";
    -- convert range of switches to data element
end loop;